import mips32::*;
class scoreboard;
    


endclass