class test;
    env en;
    
    function new();
        en = new;
    endfunction

    task execute();
        en.execute();
    endtask
endclass